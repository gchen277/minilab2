`default_nettype none

module convolution #(
    parameter int N = 3,
    parameter int DATA_WIDTH = 12,
)(
    input  logic i_clk,
    input  logic i_rst_n,

    /* Convolution stuff */
    input  logic i_val_valid,
    input  logic [DATA_WIDTH-1:0] i_val,
    output logic o_val_valid,
    output logic [DATA_WIDTH-1+3:0] o_val
);

    int KERNEL[N][N] = {
        {-1, 0, 1},
        {-2, 0, 2},
        {-1, 0, 1}
    };

    typedef packed struct {
        logic valid,
        logic [DATA_WIDTH-1:0] value
    } value_t;

    value_t [DATA_WIDTH-1:0] _internal_grid[N][N];

    /* Shift each row down one */
    always_ff @(posedge i_clk, negedge i_rst_n) begin
        foreach (_internal_grid[i]) begin
            for (int j = 1; j < N; j++) begin
                _internal_grid[i] <= _internal_grid[i+1];
            end
        end
    end
    
    genvar i;
    generate
        for (i = 0; i < N; i++) begin
            Line_Buffer1 line_inst (
                .clken(i_val_valid),
                .clock(i_clk),
                .shiftin((i == 0) ? {i_val_valid, i_val} : _internal_grid[i-1][N-1]),
                .shiftout(_internal_grid[i][0])
            );
        end
    endgenerate

    always_comb begin
        o_val = 0;

        /* Perform convolution */
        foreach (_internal_grid[i]) begin
            foreach (_internal_grid[i][j]) begin
                o_val += _internal_grid[i][j].value * KERNEL[i][j];
            end
        end

        /* Take absolute value */
        o_val = (o_val < 0) ? -o_val : o_val;
        o_val_valid = _internal_grid[N-1][N-1].valid;
    end

endmodule


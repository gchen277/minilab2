// megafunction wizard: %Shift register (RAM-based)%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: Line_Buffer2.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 25.1std.0 Build 1129 10/21/2025 SC Lite Edition
// ************************************************************

//Copyright (C) 2025  Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and any partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus Prime License Agreement,
//the Altera IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Altera and sold by Altera or its authorized distributors.  Please
//refer to the Altera Software License Subscription Agreements 
//on the Quartus Prime software download page.

module Line_Buffer2 (
	clken,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps1x);

	input	  clken;
	input	  clock;
	input	[12:0]  shiftin;
	output	[12:0]  shiftout;
	output	[12:0]  taps0x;
	output	[12:0]  taps1x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clken;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "1"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "2"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "3"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "640"
// Retrieval info: PRIVATE: WIDTH NUMERIC "13"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=AUTO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "2"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "640"
// Retrieval info: CONSTANT: WIDTH NUMERIC "13"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC "clken"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 13 0 INPUT NODEFVAL "shiftin[12..0]"
// Retrieval info: USED_PORT: shiftout 0 0 13 0 OUTPUT NODEFVAL "shiftout[12..0]"
// Retrieval info: USED_PORT: taps0x 0 0 13 0 OUTPUT NODEFVAL "taps0x[12..0]"
// Retrieval info: USED_PORT: taps1x 0 0 13 0 OUTPUT NODEFVAL "taps1x[12..0]"
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 13 0 shiftin 0 0 13 0
// Retrieval info: CONNECT: shiftout 0 0 13 0 @shiftout 0 0 13 0
// Retrieval info: CONNECT: taps0x 0 0 13 0 @taps 0 0 13 0
// Retrieval info: CONNECT: taps1x 0 0 13 0 @taps 0 0 13 13
// Retrieval info: GEN_FILE: TYPE_NORMAL Line_Buffer2.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Line_Buffer2.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Line_Buffer2.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Line_Buffer2.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Line_Buffer2_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Line_Buffer2_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
